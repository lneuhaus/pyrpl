/*
###############################################################################
#    pyrpl - DSP servo controller for quantum optics with the RedPitaya
#    Copyright (C) 2014-2016  Leonhard Neuhaus  (neuhaus@spectro.jussieu.fr)
#
#    This program is free software: you can redistribute it and/or modify
#    it under the terms of the GNU General Public License as published by
#    the Free Software Foundation, either version 3 of the License, or
#    (at your option) any later version.
#
#    This program is distributed in the hope that it will be useful,
#    but WITHOUT ANY WARRANTY; without even the implied warranty of
#    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
#    GNU General Public License for more details.
#
#    You should have received a copy of the GNU General Public License
#    along with this program.  If not, see <http://www.gnu.org/licenses/>.
############################################################################### 
*/
/***********************************************************
DSP Module

This module hosts the different submodules used for digital signal processing.

1)
The first half of this file manages the connection between different submodules by
implementing a bus between them: 

connecting the output_signal of submodule i to the input_signal of submodule j is 
done by setting the register 
input_select[j] <= i;
 
Similarly, a second, possibly different output is allowed for each module: output_direct.
This output is added to the analog output 1 and/or 2 depending on the value
of the register output_select: setting the first bit enables output1, the 2nd bit enables output 2.
Example:
output_select[i] = OUT2;

By default, all routing is done as in the original redpitaya. 

2) 
The second half of this file defines the different submodules. For custom submodules, 
a good point to start is red_pitaya_pid_block.v. 

Submodule i is assigned the address space
0x40300000 + i*0x10000 + (0x0000 to 0xFFFF), that is 2**16 bytes.

Addresses 0x403z00zz where z is an arbitrary hex character are reserved to manage 
the input/output routing of the submodule and are not forwarded, and therefore 
should not be used.  
*************************************************************/


module red_pitaya_dsp #(
	parameter MODULES = 8
)
(
   // signals
   input                 clk_i           ,  //!< processing clock
   input                 rstn_i          ,  //!< processing reset - active low
   input      [ 14-1: 0] dat_a_i         ,  //!< input data CHA
   input      [ 14-1: 0] dat_b_i         ,  //!< input data CHB
   output     [ 14-1: 0] dat_a_o         ,  //!< output data CHA
   output     [ 14-1: 0] dat_b_o         ,  //!< output data CHB

   output     [ 14-1: 0] scope1_o,
   output     [ 14-1: 0] scope2_o,
   input      [ 14-1: 0] asg1_i,
   input      [ 14-1: 0] asg2_i,
   
   // system bus
   input      [ 32-1: 0] sys_addr        ,  //!< bus address
   input      [ 32-1: 0] sys_wdata       ,  //!< bus write data
   input      [  4-1: 0] sys_sel         ,  //!< bus write byte select
   input                 sys_wen         ,  //!< bus write enable
   input                 sys_ren         ,  //!< bus read enable
   output reg [ 32-1: 0] sys_rdata   ,  //!< bus read data
   output reg            sys_err         ,  //!< bus error indicator
   output reg            sys_ack            //!< bus acknowledge signal
);

localparam EXTRAMODULES = 2; //need two extra control registers for scope/asg
localparam EXTRAINPUTS = 4; //four extra input signals for dac/adc
localparam LOG_MODULES = 4;// ceil(log2(EXTRAINPUTS+EXTRAOUTPUTS+MODULES))

//Module numbers
localparam PID0  = 'd0; //formerly PID11
localparam PID1  = 'd1; //formerly PID12: input2->output1
localparam PID2  = 'd2; //formerly PID21: input1->output2
localparam PID3  = 'd3; //formerly PID22
localparam IIR   = 'd4; //IIR filter to connect in series to PID module
localparam IQ0   = 'd5; //for PDH signal generation
localparam IQ1   = 'd6; //for NA functionality
localparam IQ2   = 'd7; //for PFD error signal
//localparam CUSTOM1 = 'd8; //available slots

//EXTRAMODULE numbers
localparam ASG1   = MODULES; //scope and asg can have the same number
localparam ASG2   = MODULES+1; //because one only has outputs, the other only inputs
localparam SCOPE1 = MODULES;
localparam SCOPE2 = MODULES+1;
//EXTRAINPUT numbers
localparam ADC1  = MODULES+2;
localparam ADC2  = MODULES+3;
localparam DAC1  = MODULES+4;
localparam DAC2  = MODULES+5;

//output states
localparam BOTH = 2'b11;
localparam OUT1 = 2'b01;
localparam OUT2 = 2'b10;
localparam OFF  = 2'b00;


// the selected input signal of each module
wire [14-1:0] input_signal [MODULES+EXTRAMODULES-1:0];
  
 // the selected input signal NUMBER of each module
reg [LOG_MODULES-1:0] input_select [MODULES+EXTRAMODULES-1:0];  

// the output of each module for internal routing, including 'virtual outputs' for the EXTRAINPUTS
wire [14-1:0] output_signal [MODULES+EXTRAMODULES+EXTRAINPUTS-1:0]; 

// the output of each module that is added to the chosen DAC
wire [14-1:0] output_direct [MODULES+EXTRAMODULES-1:0];

// the channel that the module's output_direct is added to (bit0: DAC1, bit 1: DAC2) 
reg [2-1:0] output_select [MODULES+EXTRAMODULES-1:0]; 

// bus read data of individual modules (only needed for 'real' modules)
wire [ 32-1: 0] module_rdata [MODULES-1:0];  
wire            module_ack    [MODULES-1:0];


//connect scope
assign scope1_o = input_signal[SCOPE1];
assign scope2_o = input_signal[SCOPE2];

//connect asg output
assign output_signal[ASG1] = asg1_i;
assign output_signal[ASG2] = asg2_i;
assign output_direct[ASG1] = asg1_i;
assign output_direct[ASG2] = asg2_i;

//connect dac/adc to internal signals
assign output_signal[ADC1] = dat_a_i;
assign output_signal[ADC2] = dat_b_i;
assign output_signal[DAC1] = dat_a_o;
assign output_signal[DAC2] = dat_b_o;

reg  signed [   14+LOG_MODULES-1: 0] presum1; 
reg  signed [   14+LOG_MODULES-1: 0] presum2; 
reg  signed [   14+LOG_MODULES-1: 0] sum1; 
reg  signed [   14+LOG_MODULES-1: 0] sum2; 
reg  signed [   14+LOG_MODULES-1: 0] sum1a; 
reg  signed [   14+LOG_MODULES-1: 0] sum2a; 

wire dac_a_saturated; //high when dac_a is saturated
wire dac_b_saturated; //high when dac_b is saturated

integer i;
genvar j;

//select inputs
generate for (j = 0; j < MODULES+EXTRAMODULES; j = j+1)
   assign input_signal[j] = output_signal[input_select[j]];
endgenerate

//sum together the direct outputs
always @(posedge clk_i) begin
   presum1 = {(14+LOG_MODULES){1'b0}};
   presum2 = {(14+LOG_MODULES){1'b0}};
   for (i=0;i<MODULES;i=i+1) begin
      if (|(output_select[i]&DAC1))
         presum1 = presum1 + output_direct[i];
      if (|(output_select[i]&DAC2))
         presum2 = presum2 + output_direct[i];
   end
   // Some delay to leave enough time for the sum of up to 16 numbers
   sum1a <= presum1;
   sum2a <= presum2;
   sum1 <= sum1a;
   sum2 <= sum2a;
end
//saturation of outputs
red_pitaya_saturate #( 
    .BITS_IN (14+LOG_MODULES), 
    .SHIFT(0), 
    .BITS_OUT(14)
    ) dac_saturate [1:0] (
   .input_i({sum2,sum1}),
   .output_o({dat_b_o,dat_a_o}),
   .overflow ({dat_b_saturated,dac_a_saturated})
   );   

//  System bus connection
always @(posedge clk_i) begin
   if (rstn_i == 1'b0) begin
      //default settings for backwards compatibility with original code
      input_select [PID0] <= ADC1;
      output_select[PID0] <= OFF;
      
      input_select [PID1] <= ADC2;
      output_select[PID1] <= OFF;

      input_select [PID2] <= ADC1;
      output_select[PID2] <= OFF;

      input_select [PID3] <= ADC2;
      output_select[PID3] <= OFF;

      input_select [IIR] <= ADC1;
      output_select[IIR] <= OFF;

      input_select [IQ0] <= ADC1;
      output_select[IQ0] <= OFF;
      
      input_select [IQ1] <= ADC1;
      output_select[IQ1] <= OFF;

      input_select [IQ2] <= ADC1;
      output_select[IQ2] <= OFF;

      input_select [SCOPE1] <= ADC1;
      input_select [SCOPE2] <= ADC2;
      output_select[ASG1] <= OUT1;
      output_select[ASG2] <= OUT2;
   end
   else begin
      if (sys_wen) begin
         if (sys_addr[16-1:0]==16'h0)     input_select[sys_addr[16+LOG_MODULES-1:16]] <= sys_wdata[ LOG_MODULES-1:0];
         if (sys_addr[16-1:0]==16'h4)    output_select[sys_addr[16+LOG_MODULES-1:16]] <= sys_wdata[ 2-1:0];
      end
   end
end

wire sys_en;
assign sys_en = sys_wen | sys_ren;
always @(posedge clk_i)
if (rstn_i == 1'b0) begin
   sys_err <= 1'b0 ;
   sys_ack <= 1'b0 ;
end else begin
   sys_err <= 1'b0 ;
   casez (sys_addr[16-1:0])
      20'h00 : begin sys_ack <= sys_en;          sys_rdata <= {{32- LOG_MODULES{1'b0}},input_select[sys_addr[16+LOG_MODULES-1:16]]}; end 
	  20'h04 : begin sys_ack <= sys_en;          sys_rdata <= {{32- 2{1'b0}},output_select[sys_addr[16+LOG_MODULES-1:16]]}; end
	  20'h08 : begin sys_ack <= sys_en;          sys_rdata <= {{32- 2{1'b0}},dat_b_saturated,dac_a_saturated}; end
	   
     default : begin sys_ack <= module_ack[sys_addr[16+LOG_MODULES-1:16]];    sys_rdata <=  module_rdata[sys_addr[16+LOG_MODULES-1:16]]  ; end
   endcase
end


/**********************************************
 MODULE DEFINITIONS
 *********************************************/

//PID
generate for (j = 0; j < 4; j = j+1) begin
   red_pitaya_pid_block i_pid (
     // data
     .clk_i        (  clk_i          ),  // clock
     .rstn_i       (  rstn_i         ),  // reset - active low
     .dat_i        (  input_signal [j] ),  // input data
     .dat_o        (  output_direct[j]),  // output data
	 
	 //communincation with PS
	 .addr ( sys_addr[16-1:0] ),
	 .wen  ( sys_wen & (sys_addr[20-1:16]==j) ),
	 .ren  ( sys_ren & (sys_addr[20-1:16]==j) ),
	 .ack  ( module_ack[j] ),
	 .rdata (module_rdata[j]),
     .wdata (sys_wdata)
   );
   assign output_signal[j] = output_direct[j];
end
endgenerate


//IIR module 
generate for (j = 4; j < 5; j = j+1) begin
    red_pitaya_iir_block #(
        .IIRBITS(46),
        .IIRSHIFT (30),
        .IIRSTAGES (4),
        .IIRSIGNALBITS (36),
        .SIGNALBITS (14),
        .SIGNALSHIFT (0),
        .IIRCHANNEL (j)
      )
      iir
      (
	     // data
	     .clk_i        (  clk_i          ),  // clock
	     .rstn_i       (  rstn_i         ),  // reset - active low
	     .dat_i        (  input_signal [j] ),  // input data
	     .dat_o        (  output_direct[j]),  // output data

		 //communincation with PS
		 .addr ( sys_addr[16-1:0] ),
		 .wen  ( sys_wen & (sys_addr[20-1:16]==j) ),
		 .ren  ( sys_ren & (sys_addr[20-1:16]==j) ),
		 .ack  ( module_ack[j] ),
		 .rdata (module_rdata[j]),
	     .wdata (sys_wdata)
      );
	  assign output_signal[j] = output_direct[j];
end endgenerate


//IQ modules 
generate for (j = 5; j < 8; j = j+1) begin
    red_pitaya_iq_block 
      iq
      (
	     // data
	     .clk_i        (  clk_i          ),  // clock
	     .rstn_i       (  rstn_i         ),  // reset - active low
	     .dat_i        (  input_signal [j] ),  // input data
	     .dat_o        (  output_direct[j]),  // output data
		 .signal_o     (  output_signal[j]),  // output signal

		 //communincation with PS
		 .addr ( sys_addr[16-1:0] ),
		 .wen  ( sys_wen & (sys_addr[20-1:16]==j) ),
		 .ren  ( sys_ren & (sys_addr[20-1:16]==j) ),
		 .ack  ( module_ack[j] ),
		 .rdata (module_rdata[j]),
	     .wdata (sys_wdata)
      );

end endgenerate


endmodule
